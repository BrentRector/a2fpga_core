(* blackbox *)
module ssc_rom (
    input  logic         clk,
    input  logic [10:0]  addr,
    output logic [7:0]   data
);
endmodule
